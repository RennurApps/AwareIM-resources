�� sr ,org.openadaptor.dataobjects.SimpleDataObjectj��d[�/_ L typet %Lorg/openadaptor/dataobjects/SDOType;xr .org.openadaptor.dataobjects.AbstractDataObject�]��� L valuest Ljava/util/Hashtable;xpsr java.util.Hashtable�%!J� F 
loadFactorI 	thresholdxp?@     #w   /   t GNTsr java.lang.Boolean� r�՜�� Z valuexp t MajorVersionsr java.lang.Integer⠤���8 I valuexr java.lang.Number������  xp   t HSOFFLsq ~  t IServParam_FQNt >com.bas.shared.domain.configuration.elements.DomainVersionImplt HSGGsq ~  t PMinorVersionsq ~    !t LBsq ~  t HSMCQsq ~  t UPSsq ~  t Statesq ~    t 
Containersur [B���T�  xp  ��x��|����;�%ő��N�8��,�a��ly��+�3��>�Jdɖ�Y�ޅe�����l(�ʦPʆ(-{t����I���;�m�C�����Н��������{���]��E��-���6�*��b�ܮ�¯\���c�d-b���������-�����#�zK�`�<���r�%;vY�S|�eʡ�/ص�y�z5�ś{-���0>PT�8��UWN�,{֩ʵK(�Uꕃ�_�*VE��=���{z2��a�y7v��µ���`�)[ze�2�A�a�.���z�����o[*�J�r]D	��-��.<��s
�[YZ}�~9�X�F�z\���V|�j�jN�h��L�;w����%Z�ZKV ������-�JwX�t��{:��ͱɡ����b�5�z���T���dU>��Wz}����&i�m����O�S��*�R���݌��j��Y'�O�����?~�V���)�I�^9�������]֤X��C=�|��H�/,wTt�z|�`E{(�����(X#"R��
*�rx�*dِ�-�o#�����,�K�?�����Fy�žQGԔ��^���P,y:�Jد�[�弡R��o�;�)Ug�v���t�`�5X�kۻ��r�%�g9��h�d�5�u�L�y���֙��I�Pʱ�lA�����ͽ�,2�g�+Q����c�0���ȗ����7��]��؉��!�G�{�<&O~oo�bɈ*͊��_f��C�AI�Z�H5j�Fbos�t��=,"o��^�����Ʒ���ˢǧ�-��[�bˡ���MZ�S ��XV-G���=�2c��e���yjC��J�U�P@�9�VRF�y[���xñ��? ��v���e�͛�z�+fY���OZ֢�3��E�iѢl�L�3��Mu� ����_�̉��ɛ�f�z�3�Y��3�a��R��ݼԻ5~����[Ӄzo9��zkɀ�<|����i���h��ϻ��q�Cյ��VOsS���Łu���ſ��ϣ�#�����"��{��6�ǲ65p�X���x���h�mV,�<�@O�U���.�^-�,���/c�/��v��|A�l�`=k!�!,6�>�*�!8�5� B�	���C�?#�]= X	�
��Y�Cp�!X��:{Y�T6�Ֆ����zE�Z�4c����
G\V_×V�ẩ����&)`F�t�e>�6�JY� ;"<���j�N���%j�+Z�^o�<5&�|���4U�{j�w��w�+�f���
B��i�[��eI�6Ը���p��pGT��"�G؍!�n�
�-���@p�Bp'w@pwCp;�Ap�V	+R�V--_���{�_�47ѻ� i��we�NAT��̶֘�ڬ)o�l�߭l3}�j�nM����a�n��Fe���v
���:Bn?�!x��Ԩ��Q�V�Z�4�pe�
���V��]��?�m�=+y&[��B���Y�Nk�������a�k�m���&���D-����
�����<����� �9WC�1'������k ���Uރ�]n��z�	�? ��k!��+ x��!x��!� ��A�B�3���r.��Q��l��w<��\�G|�b���`  �eu�H�r��1���HBsC%_��[+o���J#|+�5����h�^i�^m�n3^�� ���c#��L�� ��L��	�4��L� �*X]dA��Zf�/�(�Q<]����!��B����A�_�:>V�V�O��
��*A`#	̙Q��ؔ�i�g�c0٫fV�Z�i6�N����}J�eOF��!l�2\7�[y)�uV�5�f9*4��j>�W�ͧ�5ԛZ�? 4���3����5�X«Y�φ#���&cg޿U愷U57���V�Vi(,o��i��z���
-���.� Z �rVA ��4j�P�V/��ڠ��b��;C���I��2�SW�aenh`�^��PJ�JV�[Wӟ��o��$�Xo�J4V�2����CRo�dC���ȗ�����4h,�ˣ:Կ. �Eְ��!�fV.}Zn�쵫VRo�bH���^a�^b
�I?L�5h�*zOG�z
'Cp�����Ww@�o\�Jf�O�5��Q���z 0*��h�
�=+�ԬGAp$0Rc�F+d�
��
M�6�J+$c�ћSV�փ!�1��{��!X��0~��� 8�3!�a���VZa�i�
��0��B����X�
�+�G�0��B��z���\�?����H�Al�7�(��J�z|�Uy�X�n[�[R2t�� J��X��c���PZ@p��q�܀f����r�Y^\&~��u0@\�����*�]��`��*yFsggDVt�Ŭ��]��0��;�)����wpw$��W)��4��m�nH��J������l�o���P���^��(<+�B��>����e+���0ƴ��
�H�m@/�
�u+�1�w�R�7B� �C }y+���0f���z90>�B�
]l+�^�0z�B��
�u+�֭�ӷ��kn��&�)��Tn�G�'�3񓈫���n�ʻ�.�6�XC�bm��Z|�|O���!��i���E�$���K#R!��[F$:��C<�bc�KW����X�W)֗!x�?��Of��9j����:Zچ�Xc�c���6�Z>;U'��߈�7*�jG6ִ�٬L��f��S�0��AP
�0h����
�[��!����̇`gv� ��V[w�`7`Hi�!��G�Q�0D��P�
CY�<�B�<�A��
��`O��`0�� ֺ+�@ �e+��0 ��
�U+V3�Tg�2V�f(��U����}��/l���A�F�E)44�}��hgl�Q��d���
c3+�ͬllc8+����0"�mX}�q��u��}�`YK�Z���4����߸�ږ5��N��d4��Ej�m�5�Ш����^6�1>��0Lm4��{�{N�)M����{�qw��3\B����ON	��*����������+���x��5��jj9=	�<\bKt�p�F0��'@�O����Bj� �P��.��>�nu�9Y�v�6ҡ��Jht��\Ƶ����Ы�ཫ�Ye�@̯8��=�i� �|,�,J  �)A �N�	���+@�`,"@����@ ~D�W(���D	`�0tt��.Sa>�S � @�Y�޿ �@�޺ �X C,����%̄``�0��z�	`؅Rh�k��_�}
�]>~�����ь���0�5x���/�_�U��&�ʻ���Ve:�33�͆Qp�aX,���^�f��C��́z��/;�P�� �`nL�	0'��I�a� �!�C��F���`��v��-��h��|a�"��m��Z(*� ��/@� #� ( FF�!�5�
h.Y��r�ߔ�`�Sk`���LhH�i�츦4�
[U�Jؒ����
��gkA+�Ye2��l��u����o����#O�,�&k�y��X���Au�:���W���e���kcP���9:���b����(<_���VÍ��f�ot&g��x��n`jA��� C-&�	B �iX���	�c�KQz�+�0 `@.\v:-���"�i�__�n���!�����C8��a�:�td�s��M��՘X�K��6W-�*���6�ҭ���������:a�=��8�N�!-��GzqT�IRgjbM�������p+j�����X���:o�Z�#��3��ٽ��=�1��$� ��O��C��[]8���v1#���YV}F<�f`xx�; ��_�	3<�}�D�' �A�э�,v��B����]c�G�i*�϶u����������U�c�_m�\e|�rU��a���0]F���ˁ�� �M����n
�a�>^a��oU����ޤj	KV�)����� ,i�Jv� cUƪ§|�ŷ$�Q*���y��ԏ�����.�4��&g����Z��6]���{F�.L� ��D�["�D��Y���P�&�rդ��#�~�}H�+3hlX
�YF�b&��a�S��ZV�7I��t\eFF�~�͠��x�źv��D�CKc�ba�!B�"�D�ߋ3�"��x8Ի��Ⱥ�ƃ��q
V7q*���a_������MJ�V��%�ٕJ�<���qͮ��"�D
��`.$�������e��l�ꂇoI�������i�>��Хk���ǰ����G`�z&�歯F_��δ�]���0Va�.�]���GF�"���} �J)U�1��0�a�/��S��3C�b��lD�D�u�&��V����l���ņ!�kC�����m�z�X�ȯ.U�4�uiޚ�ԫW�wDo��1b���}6[K]K��}�B�C"���O[u��
��r��pn�:�Z�?�(������ZXf9�۠$aY�8	�B�D�"�*�hP�Ѡ%'��>���"�D����a�V���TD�g�l({̩�c·KX�" ��w7A�l�ㄥ=k�9��jX�%����eƨ"��� ��;X����=q)P�"�$���	�8f��`F�Y��"��Ey�0a)@.6�ND(����mC#|	��2_�HEf�a�/��G��$"��E��a��p'B�[��<`�!��@ W"4C�Z�|Y��0F��E`#-h#�u�S+�T�Q�p�fj��
�f��idՐU+Vs���bd{c;b;b;b�fXS+St93�kau�yGٚ�j6m��@[��2������Is�����Ā��$�n�X���Z�.��lU��<_�=b_���2[�����Sw_o(1��hq��ͽ��~n��x6)m�?��?�� $#g"TQ���A<�O�6��􅷨�v�O�n撉��Ͳk�+j���|E"�ğ@����R�r(���S���' 8;ğjr�w��g��s�*|�����֚6��|.���E�"�S�`�Ef��Z�`�E����%R��3�&c>�����˽f��i0�k���r�Z���l-+|�����x]�Yz�����1����_Gq5+5�ZYi�v�:� �-M��sh�A�n݅q��>�s ���h�D����&��&h{�ìj��L�b �)���Xfr�z�Lh?L�.�4+�"�__̆�|��ќ�$��j� �Y�=�|&|�Wu��<nٖ��[�ڑQ[�в]�̣V��\~��g�so������;�x1VUW���vM�wFt�_\&	��$���/��'½�DA�tr$��x���b��m��6�i3k���5@�&�P]�3XC�ٛ6pؠ�c�~��O�h�j`�.��@�Z��0�_A �:X	3�0�.�d��a�-s�uiRW��gt�ͯ��Y߀�/60�:���B�8tf��L[!�c����
�r�5巩�~ۦhT�6��%�۵L�����>>�gX��U�Dg�N�ǐ��k`�����BǗ!�2��?8h����V�_m�pz�e��㬄k�t�H9ܮC|�n�e��Y۠gm�βmO*�EjV(� �ˇmQ�h}�����xA�*¤��9H\&3Ȓw�%����a��ܻ�g���4L�xk`xf��/L��`�bcj�����`b�!�:T6/0L�A̶�m���z8�]�j�4C�G���Y%��*n]4�A n��qZ`�� E�6,?j��D);�rm0ʵ���#Z�l>n)}À�7�GC[����.��]�9�DX�&�Z4�t��[���~��p�+6l�"��9D�]�tBDX�Ǻ"�=�03!�̄"L@���?�`�j��H�y8Bl���+El�S�DX:g�1����f�6|��`"�_m����8[l�ְ���VL+Ռ�r70�@�4����^ؐ�;"�X� x�abL�=i�(�,g^&h�g!�-�"��a*Mdp��0�&�D[��z~_l�+�#D��x����!�l�x�������a��~�Wo��UwE0"��za��P������̡������
ԉeW����*�᚝���=���|5gw��GLG�wG��p�_��P��>i������!R,9z�K������0��'�cM�qj�1��Ö�6u��v���W����>v��7Y���:l���Q�ΥQ��� �k\�&1���0���	[\��/�c*�r��}��C�����91���hi�l��.o�ߪ*r��{{��_wʾ�[���=YMM�PN����Gl[`QFtb�v7��1����0��(��!s�L���(Ae��oҧ��~������-��m�=�ޕta�j���^Y��SYW3�������@|mU���$^m�o��v[��W����
����E���?��
��E/-x4Q|[4Q@�{r1U���: ժ^5$��Ʃ5�������YU,��V�e�����lyZ~��+��l�
)������]�|�5�Q�B��u��V�cψ
�=���ş�� w�n�Ң��$T.!$������1H�]K�@("�P�;4u4V��jh=^�H��Yץ�٬���x�z�dd�qG��Fƒ�Ɔ�&�{l&�d�j�qE����;��O���:W��.ۛ��'�o���_�=`��ў3�L5s"���{Vt����3x���.�z����g���"M� ֆTUza�$,Md�_670�W��_�hkRM���B����-E�>����!T{y�y���A9��������e��Xm�+j�M�bU��.%��i|d5�Z��e��V�]����߅�`-�Z��,i|Y��,�	��*_G�<������܊���鰺\g�c	:��B�Y�<H0��-�"����o#��F�э�i,5	��,�`��]^	F�$�H�,	��H�0���*��Lߙ��%�)���4	)�`���	z��9�87QT�KKl��g�������gׯ�?0\�h�~��P����y��D3(c�ẁ��=�W!�����2\?o��5��c����k6	��t��pmX]p�	�f�[l� %�`:��߶��b�^�b:�a�c	��l�9��o��z,��:/lS�}�y�`��sݶO��%�uf���~	�<�KEjAf�Ԕ�
u$��Ғ�!� 1��Qw��Bj@F%��ԊKUH�T��&�
�:��a,1�#"E�21�����$`I�8@��� A;/�WH�e<�o�9��Gm��� Z��J�趁.8VLQG[l�V;�x{}A���j���a�1�t^2͖���~]wG�ۻC���G\���U��lQ��ȶ�T��!㔂(�ԍ�I಑@"�ӒB(�	̚�S�z1���Q�"S:��1�������6l7r{����ymH�����=���^��6�g�+s	��fH�W�5[R������_��_�݊�������"�Jϟ��H'a�%�fI���z���D�)�;�HԲ��NƜK'�Τ��t�ͨ�D́�z����R8J�!���%�:�Hg����I�j�7SP���7疛@�_��o7(�2�Z:���+x��
A=h��A���������q�:(?ҥ��;G�xq��%�-"]��H?����Ө�~ȳ�ڶ��%��� �ڤKQ���X�y�T�BT�t1��c,�T�kU�1>88,�F�Ar��Y�/mU�ۦ�A����^��H����0��p}���߰��#����5�u��Lg�Y)��u��.�Yf�d���1��D-P�/�F�B���6�]�
�!�}ìu��S	�����]���x7���?�`�뤱���%�{E�`b@b=���g%�� �=�Y��C!%��3��P0�O1��1Xu�ao�!���M+�w��Y��|����4Y��+t��7�d�lX�)�i���%���/�t7�oGzӗ�B���	�Q�>�W��t.݃uE��)'U����{Es���_��2E��X~��i���|��b��ec�Xx�2J�M�_�Kf;/�U�:a�_���J�e��Z����7�d���A����@G���k>ơ��#u��cp�x]!|XW^��"?�_>�{�����E�G��g�Ǟ�/_�.��U�۟tI�ʿ��:���ŷu��Մ#�*��_�@׼�/�ޯ垑|�e;����Y�*�A�_p�ڼc5��kt_��}���MZU�1�o_��%���C���vm�I����H��0���1��}Qg;a�3*Po;���.2��{a�?��f�y��������;j<cW�e�nX*�0t��mgR��y?��ĶK�i� 	�Y݋�,����	�W���2)�6K��K4���Lݟfi�a:���Щ�?V�f]�U�9�8�u���~Ϗ=��H2θs`&��3r;�@�����:x~�a��$orGg�G�#����1x��ar4�+���ݱLEF�+���J<W�ar�T�+nX�]Q�2Ee<S�0�ʬ����$�����3�1L�2�{`*�f�๱���ͩ�i��8�����v�fV!9���<_���+���v��@�Km[;d���Tފ�[�0y��n�(r�;"+�?ؕRٚ:x����֤��3w��]���Ƀ�*g�\e.	���+z_�d(s�9��PFC�+�?2��@O���E�݄IM��g�#��7������>�/�{���s1���Po�y(�}ԅ}g�ھ;�o�sj_�y��ڰW��컢��P��]�T��G3re.%�+������X��J2�0ᕜ�J&�+9a��ɶ���OØ�g����0���Po��Q����(��TL�~&��~2��~
j�~��~"j�~,��~������v��+.�$����o¶O����v���mg6���	�>���y���&�dufso����"J`ua������������y���ڰ��z��5nuiK���hl;�#��o¶O���	��?f�;a��}0&�Pg��1����7�.(�c_ԅc7�ڱ7���s����������X�wT�.�c�8v�m����>�xm{l�n�����dº���u��ʤ�u?�w��19~�:s���w��zs��8�E]8NE�gc���0��31���P�3PO��Q㎓Q��ӰT'�;Đ�X�$t�Feoo���nrG�����>��Ȅ�m�1Ḧ���g$�7�����)&��Sb��s��wķ�=�S3K�y�h�5��ʱ�lK}"ǻ��l�Y�_;�;`����5�o���%���i3�T;����Њ5|�a�C+>���XEaQ��	��Z����M�o\ar�a�=G�/���A�V�9�o�g�{K7m��w���20B�:(�=(���k�6�;�aNo�V��� �tP���:�ƘS',��[��a��/1&�ר3��{�Ǩ7Ǉ(��+ԅ�(��L��������9j��)���	j��wԥ�X*��L���X�n��p�4��nV�,�*ܜ	��*�l'�8�p�ǭ���pH�����'CF�Wl'3�؁��5�  o�6�8`w���8�������[�O����v0Uވq��m����s�BgK������fsl�t���[��%*փe�Q�ب��h&��˄1�|~���:�l~��}����#�[��t��E�ɚ:�:� W��$9`Ӑ�]9`ە��nAl�r�fs�u�:`wy��at�v/l�r���z=a���+�I&�Dp�v�2�� ��=vp4������9`s���9��6��o��i��� ���kta������t[�$|)3�؋�(��N����k��>5��T��ێ�q�G���2������#�{��������1���pL���:���f/ƔF�ev`�3�Qo�2J�ه����ԙ!L?3�9���<fQ��S��xf�2s=�Jf�h�������}�}¶���m�Ll��[�?�1�)�	�Y�ݘ���Qo������.2@�3��3�9���1��F�è�̇P���.3�Rɼwb{�y�5���j���&I�}� ��DO�����ڐ4����m��I*������Je2�-���KS)'#��9�6�r2�}���ߤRNF��r�x*�dĻz!'/�RN����{x!'�RNF�mr�e*�d�[u��nK���x�.�dʈr�@�����,c�u
�~��g݁1e�u�u�>��[ֵ(A֝���Q��1���0�Y�b�nCmd݂zʺ5�u=�2�&,���&��N��L�-�3���m'��Ɵ��1eOB�e[0��6�[�%�v�.�%�:;���Ŝfgb��P��S�5�-�.�3�T������]/��mOu����õ�m{�
�?�cʖQg�+1�ه�޲W������P��u�~v'�4��c�������C�x��e��X*٫'��N�v��}¶O���l��o1��{Pg�7b�oE�e߄dߍ�Ⱦ�����}/�4�ט��P�w����@�g߂�̾K%����)gۣ{c'v�N�vS�>�I۞c��s\S��Y�����D��d�9y���,�:g2����9͙�y��Em�8QO99���2'K%�n�;W�/��;.Ұq\�~ھ�v��|H�q��03�8�/�����ŧ]�/��1�nF�3_ə���`�9�͊��|�͐-�1%�b��~�5�tLo�`O�	퉎EG�0��`�!e��>�J��n_�}�v��>�6�ɁsB,��A�߇�~�y[�p��^�ŒU[�T�lhp�-��q6\�bq�&���	�g+ϼ�!݋�H�u��j�e�����+��e�KwS��^�����Z��a�$���K�ٺ�?��>W�|��[ȉS`w�ٚ B�vH������eA7},T�~��E5�^{(,�=6O�X������;�y<��ս�Olw�Э�&�w�3�`��*��u���A�bۮ�;á��x��}u/����r�@���c�AN��1��w)��G�M��G���t���kt��Nj��B�Хq�N�u:U�X�=w��~��_�S��:m����B��qo��,�{d�6|)�h�D���?����C�����ifa�l|��ޣoT�z�q:�a��}�0>K7jɬqK���b3��=�f:x�w��~��^�{��7y&M\�Ow����}a��}�{�����wG�j�#���T�`�ҽؽ��n���#��nx�]}��P���?�������~9��>� w)c�t��'x���B�gw{�"��|�����R���l��{~�O���[h�h�m���q�T{r1� ��=���C��/,+�ᠻt��FwD�����׾�+�v���گԽs,�ݥ�7��&���n��w��Q�[����B5�K��l3\.c"��W�i?�+d�5=�oG#��;����F�����+�k��K�g�XjT�_�S���Ҡ�G.���;��r��-�	b����C��߾A�X��EMm?w�/��?o�be�ܖ�*ň[g0�[�v���U�Nl�����&��,E��ڪO6��q��8�ʨSI�>q�^g�������F%5Aůl��9Ȱk��2���Y��oC"ձ#?x?���Y'�8�JjlR�W,٭rW���>�*�o���b��|���T���m��?
.�)�Um���,Q�;V�"�)���&�_�6�V�}���t���V��MjQ���J��MV+�-HwO�C�P#�ǩ#1FҤ��#�0�_�Q�H�b-�5��tT�rqSܽr�_r
jY�2�t�G`I���8%�$�&K�_U��CJ�I`�s�LS	������|�]���;�Jw:4%Nۨ�ΙOE7�꜂E�ʒ�k�+�Gg6��3u��t2��/8?'[g��!n�:�+��^*PM��Uelq�{��3�߮T~;Q����[r�����"��������ݧf{{MܧU�޵˫�Abq��X2[�!EnW��X�ʶ�m<Օ����D�*���}(Os��=kj�Ofofg��J_-G��~�������C�H�Y�������Ğu�
�VY�|G%�Z�� 0cF��{����Fk[��j�=�QV�h3d��\3�|x@��(�	kĜ��	+Ȝ��q�D��xq�Z2'���&����NHԹ�U��zUŜ";]-~{�B�t���A��·���!��K�6�2"���jJ�� WͼZ}�ձ�Z7e�pnP��(P���V��vd%�����1�]��R��kA��f�K~uljfo�1rpb'�R����������:����ks�o��_ol����2:�T�{|��V�Ԓ&���(�!�\Z�~VE�E$��a�$��)�2�m�+��0X�`�[w[K�İ#�m5����EU����F���M�U���j�#z�b����d���ṃ��5�FȜۍ1�U㙂az�	՜ר�m�AfV�=���3����{|�����~���s�9~i��������uF���C4��f��&�P��R���9��U��1��m��|{�C���J`��	��8Q�YS}y�Q�
�<���Ɛ���9ՠO�1��s��
�Θn����e�K��Zk#]����f�-[�!����{]퉫7��U���e��2������^�Q��9|���+���	g ;���|6
��c�o���W�%����
�>�Xlbe}}�}3����;?��3���)T��~%��03pr�����:����f#YΧ�N:�D#�����dX'�ŒNX;鄓��p�R��\,�tތL9���Ö�pr��3$�	�ֲ5AΟC 7����	G�:_Ĝ8���㛜�#u>���	�-9�]��X7�p�/3D�� ��F�?C '29�:�|k��y`���uB'��tQ'�=���a%i�����p����5XX�XF9j�/�?��w�M�#��F��#�a����s���,���e+*�K����I���O��0nc}F��7.ftr�G�e�%��e���,�6>E5�:���STo��O%EI^�]�QROJ��)�xՎU�'GI�	(i_NI�/v��l�u�	�hi*�6�r�/���G�#::,�t�X��wu�3�8z
$��`*�IZ��&:�����t,�$�3;TI�k3���h)�����Q�߱(���$)i}J��SR�{׷�P���(���T9����I��P%e�~��>��5Շ�r�=��O%Me�&��mH�ҽ��J7Ɠ��j�	M�L��2�Ll���2o��<I#��O�g�D�uJ�d�%�#�V��
c�c-�ɵQ1�2�I�5�� Wi(ܓ��RF{KW �q"�r,���c�/jdq���
�����ZX����Eh�Ѫ�~�1L��4Ǫ�z���j�ܰy��>�66�s�P����d���U��jx�+�+	���h�>��Jl	�>Α�99���dF�oK�?^}�0�'w��C��;-�oh���	Ŧq�4�'��&��V�0�oq�i���m�lh��N�qۮJ[�G?��$�_�L��-�Z
��L���Kn��� ��A���ښ��V,V�G#�Ƣ#�A&�ra]A�*�5w9�/�S΅�sA�+P��V�gn3��"��knj%�	��Ŝ��ꂩQ���& DÚ"�DBT��A�<0�O��Z����1��$���
�I+��(U����a��ok6��4��ߐ*���*kbhC4D�*��!��ON.t�rף���vɅNi.�7\����ǚ�E:3-!P����
H��*i=�`��GS�f�hոC^Z�_sm?|�ַN6T�\Xn��I��]pk	��n��-�*���֥�V��P��c���3H�1�\��s.|�9�$�].�$ra�[.|�:f�rOArO�\��ƴx�B�ss�g2�-xZ���g�sa�{���(\k��1��K�!�'�;��5C�c�����u�u�j��?�:����TGFu��TG���d�A�!#-���P/ӮO6ԵSǩ��@u�N��{��(�Rݻ����$�mT�wS�YqW4x��� �δ$�1"�q"�a"�!"�Q"�wD�#iC���'�"��"�e�E"�Y"�y�%"�OD�s�B��iI��D�GD��D�{D�D�_�����o'��ω���_��"Q�!� �"��%��M��*����Ov��'�$�3Q��Lmr�59%���.�O��N��|x�,c:&0y&�2�25�ş<�<E�\���\�*�_����F��N��B��L�/$�w%�+҆xm�z҈�_Eb@�L�H��G��O�D�W�S��WӒx/�F�7�MD|+�B�/K�I>��2�q�N����É��D�:"����a�LK�7��0�G���"^I��'����O%1N �O&�O$��O:����O"�O!�K��%����?&�B�_H�_�6��(��_E�_Gb�������%�3"��D����k���S�x!-�����������57�"��iC���'�"�i�	"�I"��D��D��D�������R�x�	iI�D��D����W��׉�׈����/'����'��I�L�@�D��������0E�����Ļ|�%��G��SsY���P"�%m��W҉we�î|Õ�	��P�d̔+�wMB�\.�53�r�
�%�s���(�k6��r��(����/K�]3�O|�����ߋ�߃�_H��N��I��M��*ğ���/!���j"�C���5D|m��[�,��kH��D�*"~�Jķ�+���D��H|ܧH
�i$v�o��d�P��g���ÓW^�X���y�F��Շ2�z15��r��(�+b�E�g��X=�X�[���Ī�X�@�n!V�$VכZg&��,3Þ��bҀ_�.}�:|�u4�b�|p�:6+׀%�Z���:��_��Eܑ�p�/�۩��V��:��`Z���K�!qʮ㸊%�!��0��6�`.�x�ôe����&�1��׮�3�lU�u`���Y��p�e�u
��:�09��b%�m]��|��Q2�9�ę���P.�"�:��ش�5�����]f׉�-�e�^�����SP]j�	�rm�W\Wab�+)ڟ�<�� �Q[��G�gX�^�ҿ5�X+�����$6�U�_2jc��ͪ��;��#j*��;�n��t��8�"��h�@��[x��-39.w����`P��J���B?
;���N&��}��#�ƽ���,��M�q>s��9�[`��/uװ竲=��*Bу��b���:r�L�3�YP@7;��$'"�*�[�a>]pj�/�i]�u��u3m�n�6�'�_���U�[��-Vh�ä��9ڄ/�8��[ʫZ���P��p}��x�"�����O��4f=d��
��ME���7݇z�A�9
�ڇ�u}���>��N�V9ҫZ9�F8a��ϷZJ^C�˴�;ǭK����'P��,]o"�?��\G����u}�4�^�ru��ֱ��ǲu��t
�����`f�Q��q��b`]w"7��!��ɮ�mן�,�e��V<���3���`��Ul�.����zu���L�C\��e��k�	�א(,�e��+�Y�s��jLc��l�,�>ke�`k[vNo�a��w�{�͘�Eϳ�+y�X����Ij���24LF�L�V��N�N�B����G��3M���؞��~y��b���;ۑ`�M��I%�O%V �L��$gX����t��AټY5�H�A���؊{��{eE��L�G׶���5�Q]�/�U@[�W���C=��>x�A"�Y�<�sص<�/��0��|*�9�]�ά�;=�&���*��Ư�J"��n�:&H��Dx5iu1~ K�ό���<�g��z�H^+�E���h$5��H��+Zy�d��k.yG��1:A$�P�_;�o��0�	"��3��]�㓖C<��G3��i:e;.����P�дhۭ}�����0�C�6ߺ ���V[]U��ɨ���q5ѧ��o;��{�Sã7� j�Y�7[�uu:z���/.����<��1�_�˃>d�������A/;�U]%Fu����TgRCue� ��:�V��[mq�8�����[�A1T-�wXx��·�<3:X� �կ� �����	��`J.��y0ñE�u���y�<�fQ�c�RC�/�}�x�偛/�m��j�|��E�w
V�< (��y�5���:�л�c���y��4h/�j1sy0�cm�^Xm��x�<�@���x3���c��~l�S�)�Տѝ'���1��^�\k����>���Oճ�$�o�<��@�d�}��5���u9�Y�*G`%ҏ����α�G݌��݅yͻ��[��(��̗�T�"�Fx�4�f_ha%�%�����m�����Oey���t�ũ���?)&��<)/v���d�׏�Iy��5���˄�L�C�qBr
��5��G&�����B|b'��a��9�?n�'GC��A�����Ґ�Kl�Y�ڟ�Ѫ�G�%����Ҕܱ�i�(k���or�J�C��*��QT��u\/}Pdx�=e��`j�PZ��޷�D)>�U|a%R��7Fn����o�V�Mp�Ք�c�5��99\%�)ݼ����5��hH;t=���ǣ럈��N�����9�?�~��ב�/�D�i�qZ�r�����h���O�C���!�U�GN���8�����;TKR���$GI�	(�Y^I�U��
�MJ}�f�;����(�횙����N�_��-&6�+�v�7�}	�"`~�>�����3�h�6_�W�1���D��8E�3G���s�t%�I��r�:������|�V�h�*�H���0��X�p�3���|��/������/�����܄���PZ�e��:�W��=���������	����9H�[���>� ��h���&�`2T<?�;��=�RF�'q�G�����T�K���CP��Z�1�S˯G���P��%�'1�J�N�>�|/>����_����L巡��+P���(B�����婲7-O���!�D����&�D�z"~C�/'���D�1$�V"~$����B�E�M�oN��r�y��D����3��3��s������ӆ�S�O��D�U$��D�v"�
"�"�2"�J"��D���B|Z���;#+3K�]򉿇���x���������������_���'��DĿL�?G�?KĿH�?OĿ�6�?�|�� ��Fb�CĿOĿKĿIĿMĿG����+E�O���%��E�I�A�C�E��6��t�
���lcj&05E�j�LMQ��
6Ձ"L���N��
�iyb����ԙ(��"�qj!�6��:%�:=]����4���$�"~"~'"~.?��ߙ�ߕ���"�O�NK�"�&����������$��%D�2���o&���z"�"���o!◦
�iI�:"����!8�#���G��k�O�"^!1BD|���%�D|���#�#D|O��GZ2,"<B��-�ğM�_Db�G�_@ğOğC�����1!n�����$�WD�5D��D�ψ�_�?'��6�oO>��%1� ��"��$�o%�o'�M�����-E��b~Df��"�I"�1"�Q"��D��D�iC���'�"�/$Ɵ��?��/�/���/�����ͩ� ��I�H�@�L�D��=m�?���XH���G���������_"�;"��!~�;�H|��/�CI
�(cA�V0�*�����I'�`:_Fb�`�Q��Y���`&
V�F
J1�3R���Ғ�=�����݈��D�D��D���!~�� _KbT��D| 0�!�k���R���Ӓ��D�*"�Kķ�+��6"~y�ߜ|� ��$F�E��D���o'�;��n"~]��lZ���?���H���[��MD��!>�|�O ��$1N!�O'�O%�O$�O&�O#�� �O�͞>��G~F���8V���8~_�(���[c�k��l�:��b�+cbR�?1~� .E�}$����kt����gG��ZK��)����%�e
��m�w&y�ύ�Ɏqy\5����*�k)���Ӳk�q0��!�/n��FO&�s���B��@�2�S
�	����辄��Y���K���Y�����U��ΐY狰e�&'�|��{��X�X�*%�_ׯp%���J�pr��j��I�Z�Q8�1?6�����N8�a]q����_X�!����/�I���TG���g��kA����D�&f<
|�І�Z1�Bq��ˤ���T|�W}����ܜ_��/N�����T*�T*��T&�~s�bɨa�%ѕF,�dlЇ���}�A��q�/��t����#r��KVj�r��=��
�¥g��/-+u��֫Z��b���'Z���{��Y�迍�@���;��
�P����6d�J�~�N_ "���n_�K}��?���|y������R�`	�����-kۂŐ�8�P,6���ϓ��F���I�C�}�/��M���as���%Ǔ�ޖ�C����P�(c�
L�p�U�
%*\�.ޖB�v�$oKa>\�Cbtc�P�B?f�PF��P���(Ba 3[ؙ"�Ŝ�\'Px4����B�o#�$�J�7&��S��sI�3�����3��S��Ӊ����s��ӆ�/�c��	��}������߱��#�_��^��^F�^1�#����^n��J^?�^��kFZZ�Ri�N�uE{ۨ����'TԎ�Zu<������X:'��/>9F���G	��	�G��L��@�fn�BX�;�[����|H�������N���ՉP:đ��w.IV+��*����|��耍�Y�1���"�q�%ac�1*�a<�	�{]�WN�w�C9A2ƥ(;(*�9����C������R����Р�+E�1��B��h��	����h�T��9i�ʩ$v��(���3q���	�f�*���=8�����h>_@I��PƢNL�h=�Uԍ��ŃSԮ]'ɃS���E�H�͘@ё(J��TQ?�_�	+ڊ"��-ژ">�"[Z6:��4"�,"�"�̴!�����ĸ���������		9%q�_�YZ+=3#S���	�F�o���I������������{�������{Rgp����/zD�Nl��4�R�&V�E����*�����^��H��m*�w�<ޢh���=���Wi����	}�k���C���R����^��ė��	�ڋ��!|�p����ڷRY|�q�jol��D0M�w˧���ϧ����i3�i%#r�۫�YJ��8J�t�K	�����@��u����8Դ'��Y�P5٪U%%GG��\����Z��]�_G���D����U��F��~����>����I�`�G���e۱5nu�j��j�Q�T��5��j��J#�(�V�&���$�V��c��[�qAc���[�c������$u�'P���#�}p�ar4��Z&�NC�wh�hl���hI�N��ꑱ��cf��f�{���)��9�(9:��_ۦ}��h�W@G�'GG	|XyڿSIG�ʕ��!9Jꉿ�Mw�Re�l	�����w��'��8]R,�Œ�[kjkZk�<5k�V��P�k�\�9hYY�(+�3�����V���x�r�ũ�K�`v|�L��l���d�/ �K��T����A�G27o���{Ȍ���Y�^Z� V'ӿ��Yޠ�^M;ؿ�Q���H`)�􍼚v��#�J�X~*jڅ�*�Ա�v�La��c�������䀵����s�X�kL�ԫ$GK��~��ZڱV*cu��	h�>^K�xiilWĴ��������/`bӟ�h�??����I7�|i��c��`��T�SI��J⍉������o��JI|-����x>_<%)��2�1��r���%*.K����3��$�E-�����!1a�{�(�{`����Ż�`�{��{cf�wK����7�%�K��z"�����uD|_�6�k'��eD�c9���_Aķ�mD�J"~5�M���qŴ�����Ӟ�b�SVL{ʊiOYq��)+N���b�SVL{ʊiOY1�)+�=eŴ�����Ӟ�b�SV�*{ʦ홖�Ӟ�b�SVL{ʊiOY1�)+�=e�i���8�{ʊiOY�v���Ӟ�b�SVL{ʊiOY1�)+�=eũ��l�UiI<�)+�=eŴ�����Ӟ�b�SV�6{ʊ�������Ӟ�b�SVL{ʊiOY1�)+�=e�񴧬x���E|iZ��"��G"�y"�Y"���!����"�}�-"�]"�m"�u"�M"�"�="��T!�|CX��5��9����e��Ϥ?Â��D1f�0�ve����aE�g�(،a�3;CH�;ӑ����$Ɍ�q�TLm�4�kF!J4�(]����|�ˈ�]H�yD�ND�|"����K�/ �w&����V�%���? ��%��'��#���{%��Z"���XJ�7��uD|=�@�7�KR����$�"�G�F�Jį%�'��6įJ>�~">Lb��D|��_O����G�oH�_NK�O �O$�!�&�'�%�K�L>�g������?"��"��!��#�Lğ�*�?�������%�S"��D�ψ��ӆ�+�O�MD�]$�mD��D��D��D��D�D����[R���%�O�'�!�G�?N�?J�?�6�?�|�#��Lb�DĿBĿL�?OĿH������!U�� -��;�1�7"��D�GD�D��iC���'�K"��H�o�����"�"�!��M�����:E��ޑ������gNFIff��3�0���P��9(�Lg�?Ӟt�g��3g�30���P��31S3���3I��%(�L7fv��T!���$~�_A��J��N�/$�wK�wJ>��j� "���?��ߟ�?���$�=D�)B���Ғ��D�
"~�Bķ�D�7m�oL>�?$�H�uD�Lķ�k�x�A�w�G���OMK�7�[�x�����~"~c��m�K���'��'���'���'�
�ק%������?!�/N��O>�W�7��"�#�!�N�����������E�IZ?�["�7D��D��D�=iC���'�1"��D��D��D��D������?�O����NK��"��&��BĿFĿIĿNĿ�6�k��H��� �?%��I�D�L�B�F��=E��>+�/���%JRb!���JD��Ċ�iC��N|�.)@1J\�@I>�R���*���LF�J��%S1�%�F��z�|e��md���i�	�rR2_))��J�m)�������,�q��P�.#-���<���ؓ����W�p���jv���7���F����&|����4�o����%��R�L"�*�����c�T��o���T&���I91��4����^�$D�2#���@K�S@	��D��^Kq��8����G���芾��<{8]����j�Ni�SWbC�k�*J�j4��͞�5Mm&�P�H`���>�خJ�ri%��ؗ�x�T�hN�+�*�9ͭ:x|��Ԝ��K��G�R=rԄápcd��)�#���%Orz��C���U|��¾�$̜���J^�45����lh�����j��]q4b�$����0�]'4�e�Wfe`b�D�v�4q<�iWu�T|iV�;k2�D�D.��k�x؉�a���;�9�R�D(�$'f���g�BIfyQ�Y��ڬ(׬6�h��t�D�լ]'ia���,?�с	��BQfɘ�Y>V;
6�E�Ս���.E��&����o%�$�7��D�"~�9m�'����3I�S��Ӊ�S�������ӈ�3���R���iI��D�D��D�O��ˈ�K��Kӆ��O�/���H�k������_�����7�J�K�LK� �$��!��&��'��%��K��J>�O�ϑO���O�'�$��H�?K��!U�=-�������������+m��s��;�%��	�9�)�1�O"�3"�"��B�E�H�;�w�Q��2����[B��"J䶥���t�ݹ����pO��(�;3垌��P0�T�]��u�R���Ғ�D�ND�"����O��%������'~���؛������/��g�,�t<�>�h�	�[�k��L�]C��}O|���w��{�H�c��aT�)�CG�ೀ-����j���;<�!��^�X�9��?�|ɭ���Ow���Hp������Q>��O辍����T���qQ���ڳ�+��ƛ|��zv�4�И�V��H��ZP�D�#X�X����׭O^I%�(�m��x�$s^\�r1U)�r8R�6%kQ�zRX�
3|�z��ĩ�PX����-@�.����i�q��b�г���S�M��X=�~�S�x-kK��P�'yX%�X��6�ո٬1��7Ҏ�W���L��%E��ĺ6ӆ{�_���um�|ev�u�Kb�8��mb]�� �{�ڲ�UJ�RwZd8����%�]�2ή��f/A�fעD����W:�R�N��tv+><�Pc&0{5�2{%fj�ş���
E��3;�-Ef�Ϥ%�"����&⻈�D���_�6�w$��~"�hc����H�o&�$��R���<�j�9D��D�D��D��D��D�YiC�)�'�'D�OI�ˈ�+��ˉ����K��+���D�%�B��iI��D�mD��D�D�-D�MD��iC���'�n"�w$��D�CD�D�=D�}D��D��D���B��iI��D�KD��D�3D�D�sD��iC�S�'�u"��$��D�{D�;D�D�[D��D��D���B|ZV;�"�["�"�s"�k"�K"���!���_jŇK�P�R	(u�(���R�/��`�v�43[*��*����]�S��]'��-����bb��m��t�Oi����)u��<Py�L�1���i��u�����z,�N�$����
_*��Ѻ����a�������a�X��sl���,�zqpڗ�S���OƩa��5��<��kǈ��ؽ�����JrJ)�e<���_J��q�I�x��!:�-m�44^',ũ!�*Y*
$��3SIE��p����#�=%����
��u�P=�+����3J5%x@����5�N���K��w d�.}&���қ���U��V�F9�u%ie[� K��m�&'�&�X�)�Z�������<9�J``����_�Qc<H>B�NhTT��W�h�Y��-˜Xh��/��/�M�E�e�T3�$�PIL�X8��L���E���*��ࣲC����P���(c�
L�l�U�
%*[�.S)e^�:IS)e�pY�э	�m@Q����2�/�B��֣e�lYg�L��������c���D�"~$T��1�ğBğKb�AğMğIğJğNğEğCğ�*�w�%�?%�"�/'�/#��W�W��'��k���H���[������������[���S��/Ғ������������$������H�g���������g������?�
�W�%�%��FĿCĿMĿOĿKĿ�6Ŀ�|�?!�%1� �&�$�?%�?'�"�!�?K�oNG�˳���l��<e,�0��L��܎�;҅�r!�ėO���g���@�t��3U����`��P�r�l��T!~kZ�+_A�/ ����;�;��s�O��D�A$�~D�D�b"~"�D��D��D���B��iI|���o �!⛉�F"�)m���,�W��H�É�#���k��È��D���?4uz�w��B�rm�mb3u�=�Jy+P����B��#�w�w�摖�qT'PyK�?�ޓ�["�����bǻh�-��-@�Ε�并n�b�>��{����n%�(���V�ew�%��&��;��;����
v�����;��ހ���)*�G�}���������F_�]���%��j�>E�a]�_G|9W	�T0!]쪔� �����U���ՠO3����������r�������h9{�E�����OL���*��)�u�[�m����pQ;;���_f '��]�d�Qr�u�
W��#T����CO�bݜ�ܯt�T�kz|���ېH�l^;��9��9��GkA(��[��Q�cx�vG�{{Ca%�Vv��CJ�=`U!��I�����rh�y����C�+�����ЈV̻�RoQ�`�}?f�}�j�GX�C!���=�df4D(� ���Ö���_��}q���S9���#	5��h���5?�SMIm�XR�F��R���_ᕿh�*�Y
�my��7r��e4^aиzmR��P@5~��zC�F^m�Pq(��W�8����r|��݉�R9����[�n�T�Q�|��Ƿ����@�C��'ծ����C��Ճ6���J��o���cP>#h�ՄG����ڇm����j߱�j}�=�3u���W��R�c���R$��~ΜT���j�E"�Bᄎ��t����RI��J`�ٜ}�+#��AcXFG�]F�^��X:�T*��\��ҠڱCFH�÷*?�՞J�JK,�c���CԉX*n_{�Z5�4�z�����=�6t��(��W�v����&w����+�%�VƠ\�/���<��2��G��N$�sb|&)I������Q���0���E)��6���i�0&��6�DD�����m3����9��c[
���a�p��}aR����IR�O�ݧ]'4�1�9|e��؜g1�9Ϗ��Ӝ/Y"�2�^l?���4��1�~:�u*���$�B%��跟*����KDW�ؾ�[Pmw¯�܂�X�L��o����ݨ�W�b7��a���z�9��jR|���y����(��2�qn)�6w.�5�%�;']�{͝�]'i������? 1�����35ww�(�ܽQ���bf�.J��s�%�K��C��Z"����'���%iC|U���+��5D�*"���_Aį&�%◧
�%�=D|�����D|��_O�oH������?���J�o#�$�7�[��������ͩB|_Z.�#"�L"�"�"�,"��!���1�q9����������������)i�mZ;#+3K�]򉿇���x���������������_�QZ��2��,�"�<�B��t�������>�.�&�6��W"��!����$�["�_D��D�D�7D�WD��iC��I'~����F1�e`�2Q�yv��<ş'�`�(¼,��<[�?g�t$~�|~�L�d^�8�S�Gr͛�͛�.���O>�s��
c��?���O��L��J��K��_IK�"�&�������{��Fy�q�vv���$$!��a����W�I<"�a'Q䳭 K�t� Z�0� %����u :�b�tPf��I�d�@�%��s���aپ���.�?�N~���~�ϸ��>��癆���'�\�b,� ��ׂ�E ��7���F!�)S���A�2	����� ~�i��P�/�������A�� >
�;�B�^S-�����A�5 �j��4�N��@�M ~3��*��
�����o�7��Y�LI�= �^'����
���w���o�O��@����0������?��?1�3�oJⷃ��@�� �)��?�5�џ��A�N��:�Ŀ�_��7A���A����)������� ~����{MC���'�c
l)�@�a������OA��B�23o�H�-�HK	�hG�Y&�\�R��2�,�[F�N��x?bL�,'�(��P�o�F�Y8�r�2������|���d�֪�p��N9A���|��g���=���gM�,.�bqSf'�-��	zR������2e~��n#��g�����,g�Zհ�X�
���|�c��ԣb�Zl���Z��:Ő�-w��W}��J��`G�At�K(�eY����:V���@�Y�c�e�Zَ��(W��~�:3��{�gޓb�DJ�`ˌ��F��vBKu��
�_nO���`T���fiQ��Hn'd#8��g��Йq㘹��ή�O���5�
&�&��������yy��lo��n9�
F�ґ\G�U��VW4W������[�3�(���`��*�(V��5�vO�Y�G�������y]��.��l7���2=5�\�R����LWU�g���LUKbbd]�	���QW����յ?M]E��K]9~G�"��il-�(�ᔙ����d�uPg�L��G�� �xX�XX���0���Y{R,�Hi���ޣ}򰾴:trAJ�\�\0�_�h�}�<b��w�R
o=�$�zIF����BrY�H"k�Yf߭��g�f߭�)��b�)k�bm�BYW��֕$�U$��TX�� �M��$~����@��ׂ�� ~�i��֟��A� �F���o �ׂ��A�� ��o��i�� �w�����- �v�u�i��E���?�������@�� ��]�}��(�MI�/A��@��@�� � �� �1�����?�1���σ�gA�v���o3
��MI��@��A�@�N���#��4Ŀ�?�{@��c?�������@� �� �=��ӌ�ۆSx��Ć2�
(7[1�e+$�lE�!�����J)��X�6�2�M�؎�B�Ɠ���$�m2�`;�
k�Ї�����C�65�b�)�gM����(�m&ef;��ȉ�S6;<�8>`�������ǩ����)H��A����W�`�U]�����q�+"FŐ�|�ۄ�{P�m�>�i��X㋈\mů}�#�N;í�r�Y��l�֘#2�B��[�`k�f2�><Ȕ��y���e��H�KcS�Ǵ��ˑ����~��A���E"r�P�sL�:���^����O)�r�}����4����v����ʠ��O��_�CiE�סּ�6�0yU�43��\i�e�i���U.�>n�*Wt@>nÛ;Ĝ\�������=!��7�H�]�n�<y]�ª�;�9�)^�B�B/
�s�L�a�:�A�7J��-å�P��
5��t=Yz��0]�T�m��5e��1\�!�[�{ ��%h�R��$.�[�IZ �W������'�G���8�����a�fW�e�v'S��5"�$v}�raMT��b/�[��&�3U��_�X ~�P8\�����ܵG��n?L��i�a_����w��K�����[��R�	H�;����Y*������#�u�$�z̆i�ߏ����`6bq��梧��c,���Yf 8\��^I�_��Ym�������^�vS�^�̶��r9�>�>@�ls�rh�,q����x��p��0� �{.�%�*E��q3.ܔͣ�e�I��3HƲ�)���$W����L�,ܔ��|�i�l.k�)��:�l�����+[L"��Sa��5�R��S���@�� �"��_◙����'> �#��w���_� >�A��F!ޔ���m �׀�+A��A�� ~=���4�_�?�_�!�M �� �f�%��	���l�_1%�w��� �� �[ �.��i��?����?1~��?�?�?����@���B���$�Y��?	� �π��@�Ӧ!����{��xĿ�_�/��W@�� �M��Q�_cJ�����@�� �� ~���w�����O�G �0���?�?�����@�!��Q��ߌ���Sx���>�d�����$�}Id/1����o?��O�S)�	$�}�>�ķC0�t��Qa�����~r~�l�3�Ϛ�-�v�bwRf�2$�8B�l�s��dk?m��8���=�B��>hq�r�bu-;��3=Y�$~�������_@����/��.M���7�Xe�%�_��M�������[�[&R
Ö~�}�9燚H��s�J3�4�j�z󸋁r�Z_.v��d��H입�X�f�S��@��y��\�u�WP����i/��Zu|7����+�A_���/�c�-����,Kv���N�d"ݛn�#�pNVȇSi�s9�ʼ%�&W��ȆH���6���*3TerYeV�'�=�[�2��$_D[B��4ZN�e�-�׸���R�r��!�uLIWT���h$�r�>��pꯣ�8��?J7飡�z�f���|�(�Y���N�a@E�T���϶u�	�&b�noW���߷+Ǌ\�J��U�'6�&�5�d9$��XM��O"`�:b9٪P���1�2�Vǵɱ1G[�a��a�+a��r�Ua��K$R:��*�RΏ��V�񶾴:�U!%J.�*ݯR�/;��q���4�w<C�8~�2=N�9�"�O�D�'Ͳ���e�Y��oǋ���x�2p�F�8^�B9~G�;^"����ש������QfJ�w��= �o(�_A�.�w��i����������O@��A�� �_ �? � ���(ď4#��
�,%I��IF�(��9��R{P$r�5����<�;O��S�i$��rK�;��`Ω$�s:�y�Q��7%�� ��� �Ļ@��;MC�E�� �c�?���s@�\�� �g���[LI|�o� ��{A|#�_b��O�� ^�+@���@�% ~9�_	�[A�2�o7�v4�j��G@|7����(��LC|H���C� ~#��į�W��kA�u �*��aJ��o�A�- �k �V��4�߬?���߅w��{A�V�������4
��MI��A�c �a�����?j��?�O�� Ƴ �9��?���A�� �i��XaJ�����o��7A�@���4Ŀ�?��� �^�Ŀ�w��= ~���6��Mf$�UH�]E �0�?D�����OI"W�i��Dw�]c)�k2��O�&�(�	T(�8�UJ��&�������_jN�g���I׉$���3I.�I ~�Y�wMӟx'�?b� ���.���?ė���x"{�U��Z��-Ǯ���r�:#�����UIQ\Ք���V�j��Dv�q�����U7P{,�=·=Z��y��r\5��gJ��r�
S$WW���V�p �K5o9v�每-ǊguN���-3��P���Q�P���hPDʳ���`U���u`�y`��٥^~M�$�J��[ɵ9�J�>̃�X6_R��'�ѐ�'�H)O�5$��hm�[�|:���^*XJ�ɗ�;(Tjj�r���¶zږ��<maR���LO�b��GQ�ڑ���5N9�~i���)����k?��`h�I�N�|E*/��N�A�R^K�%�4�i�M����&}��4�Yυf��,�����$I�Y$c�|ʭ���*?�$*�0ˬg���g�f=�S����H�7�(�K�P�u$~y	V�%ʛ�������)�o�� ~%���x��A|�i�_�?�a�bDA�j/��.�1��w�x�æ$�#���_��A�u�!�*����o�������- �� ~3������bⷙ������{@�V�]/���4�ߩ?���_@�G@��A�� �A�0����?d�w���߂�A�v�Ŀ ��ϛ����'�u������w��7@�[ � �m��Q��lJ����	�����@� ~?��4��֟��]1>�܅$�� ��I0�0�]��_�=:��:��gM�����=�2s�"�	G���{Z~�u���3`�Y��IHv��u&+�:�zV[ $�.��MG��wg��J��`G��{.Er�ˑ��4�q�8h�ޛ���oug��q+e��w���wg�=)�L��[f���bvTK���<���.NY�f��f��q/����3�����h\,��Q}̥����O7�'y0��"U������́GO�'N�ci��=!_��q�{�@��(�����z${cN�
�}��{/gJ��m�}{��
ܛa�;`�[`�[s�V0kO�%)�n�ʼX��
N֗V��
r�V0�_�h��q/2��{�w�$Iܯ�L�Qn�H.�$��M�Lθ_N>�49��+v��(�^Ž�
����~�s�!��Qa�7�t�;fJ�?��|�?�2}���� ��i��Xw��Q��Hb��(~<�P���$>?��KI~�c��f$�?	�� I��$#?�r�O$��H"�3�|r�P7��@� 1\ ��� �� ��= �����w��g�w�?5���}�?����?ɞ��	x������w�_8P{4�-���6�5��"$&�P��P�KP�Q���J�jBR@
�ѪpH�Bbĝ,R��H|6C*(�K�����vZ)a�MlHU�p�s�/�v�"b��5�)���Cm��XD���b���δD!�!fF���-fF�%�e������R��'J�g<�9��/ڐ򜱇+%�uF�Y��	h~#E��:=��p���
�Q�Μ��ꭻM��ג���d]^"���Ȃ�Ƞ_.g�)�a߮ ��\�O�^Y�S60�vvSdS�������R�$���u���w@ǫd��.��&g����hl�jjl���L����pF�����Q����ȫh�hcr9&=�a���(�j���2��g�Q��G�[A�]��C��g�-��K��������g��<[X��g?��]Y���@��7QE�%�ul
����n<��q��7��g䭲R'*Ÿ����׶Dͨ�T3Rӄ`��x��v�kE�X�ʲT��sN�p��XV�v��$Y�p��)�rA&l�*<�gr��'��t�w�RA�<\����rU��荥��*��5��/��߳v�"Ä1�b�L4���xJ_�<�4��.����Ӄu�6ZP���ϫ�xo#�;r��J)�"q�R_0&�,٨&1�:���c'�:�zi����$��^Z�tO�M�}z5��p�3�U�9��l&��K7��;�f�K����g���l�g��<;��g���̈)�m^וR�����O�7�>D�/K4-kU��뷶��<����^�����"�~smr�o��Q)�98�#��<���t�9Y`���!r�uQI����1���������c��/�sO��9���8DQx����a�NGg��J�P_1���s�T���`�U��Aџ>��N�(�U���5�Y�aps���_e,*����k��?Q�3��CP�7����$�(�OW5I���La㜚�rO��맵(R���M[��\z�\��~*��������'��-C�IQ�4��!BU��-����Hcm�"n�����]!7�`p���y�8�ş/`֊H�Y^e�K�W���U�5�d���?��������c�E�Q�c��I�s���dA�W����;��̰��x��nl2g<��o��;�ّ���xve@�1#ᙓ��YU���ꩢRy*H���s.��!�<�P>�E�O%��SMRy���ڵJ&I�Q"���č�}*?[�a}�g~�.��}���^��i�+GizC�O5���LM��=�;}��t�,�[�=�~_Co�)�h��o㕖D�*�g�T0����+�/T����|N���(�R��(tIS{�4\k\�ٜw��𸒭��xʿ<)�O���(�����=���,z�+��
��Ҽo�`�'̼.G6��?��fbmפ�	�DI
�ڣ�ڐ<`����Ä ���p��m�Z�k���Ts��QU�y����?��_�[�ޅ��Rx�//��vaJG$�
���s��s�)^����s���m\}C3gQ�W=g��ͮ��h�m�����%�yk��\�����y��%�V�x!-Q�RN�$E+c��e�G��XFvN�&7
�:���6D����Ґ��!�K׆�Y��^�=�EزO�<]���K�y��&�r��gm�%��U�� S~mm�D��<�����Ҩ\�|�P��.�5ae� �Lħ	|�2���@�ŧ옎_�u\s~mSsS�o&?w޹5���J���l�o�=���WQ_�����z�����r�o�Y�L��eKJ)8"�[�:N\+[0����/�
f�!>�5��&�;$)�sd��ZB�����p[��T�ST1~I ��6���Z*��L�d�Θ�T���Hxu�Ul͑:��X��Dć{;'`n'����*�;��g��o#�?�����n��-�UW*G�g��j�4�S��P��ԄV"��1��j�����0���FU�T/������kuMSUگ#�_���V���X�ZoS�wi�?F�T-�hJOc$��Ż���ޞ�6z���|����"T4g)XsmFq��Z*�x{&�|A�xC�3l 0�=��P�>X�X�؈A`B`b�R+������z�F���
G�f$�m��`A`�s0X�%$_��}���a���"�e�A&�y�>N�-�S*��o�髬#9[��(��P�>�$��"��N$��
́�f�dr7��4�Y�Z$8��R�������ȣ���D�!W�B~<.h����Ɗ�CKu��6�R��$�ì�a����>���X����tA���M�?J��j]	+�-�4!a�F_�י����[J����ϖ��򴆦��>�L��xa��ܐ����_p*��=�ZJ�
U�l�M�
lU8����p&��C���M�
);��L(�FEjH8a�b�m.�R8��.,`+S	���4��MAPݢ	M���|�z�ˁ.kz�V5��&��`K�nO��L�^�O�T��|6�vT(4�-�)��̄6$���M{C�h<����K�=_S�M�X��ٕGc	�g�*�S�yEV��Pј����)=L�7=D���.-�"�W��!�C}�*}�������~��4;Q`[�vΡ�EfoV����rV0����������ܢA�r��-U[VaC��Z�ԗ���	�CN`r�V������j����Х}�(��D�<'�ۏ�o�y�T�ի����̫P������W�@�̏W`n�ہ"�3d���(��Fv��܊�d(0�A��E*�cH�o��'0�U��� �C��5,���/�v$�p#��U�
�}�e��W].�;�GS�����	:�8�Q���q^-�>�G����6�������/7���[�2h���Nx�mTk�픤�E^�d��YO[��TE���)��4��0I���5�|	t�
t>�\K2�N����wt HSGsq ~  t HSRZsq ~  t MinorVersionsq ~    t HTRsq ~  t HTsq ~  t DomainIdsq ~   �t HSCQsq ~  t PMajorVersionsq ~     t 
DomainNamet Test1t HSCLsq ~  t Lockedt admint HSCHsq ~  xsr #org.openadaptor.dataobjects.SDOType�s��Ԭ=� Z isPrimitiveJ versionL _uidt Ljava/lang/String;xr 'org.openadaptor.dataobjects.FixedDOTypeDܤ�]ց L _checkedTypesq ~ L 
attributest Ljava/util/Vector;L attributesHashq ~ L nameq ~ :xppsr java.util.Vectorٗ}[�;� I capacityIncrementI elementCount[ elementDatat [Ljava/lang/Object;xp       !ur [Ljava.lang.Object;��X�s)l  xp   (sr (org.openadaptor.dataobjects.SDOAttributeJE+���1� L nameq ~ :L typet $Lorg/openadaptor/dataobjects/DOType;xpq ~ sq ~ 9pppt String        q ~ Gsq ~ Cq ~ 
sq ~ 9pppt Int32        q ~ Jsq ~ Cq ~ %q ~ Isq ~ Ct VersionCommentsq ~ Fsq ~ Cq ~ /q ~ Isq ~ Cq ~ q ~ Isq ~ Cq ~ +q ~ Isq ~ Cq ~ 1q ~ Fsq ~ Cq ~ q ~ Isq ~ Cq ~ 5q ~ Fsq ~ Ct BVersionq ~ Fsq ~ Cq ~ sq ~ 9pppt Boolean        q ~ Xsq ~ Ct SCHq ~ Wsq ~ Cq ~ q ~ Wsq ~ Cq ~ !q ~ Wsq ~ Cq ~ 3q ~ Wsq ~ Cq ~ 7q ~ Wsq ~ Cq ~ -q ~ Wsq ~ Cq ~ q ~ Wsq ~ Cq ~ q ~ Wsq ~ Ct Pswdq ~ Fsq ~ Ct TPq ~ Fsq ~ Cq ~ sq ~ 9pppt Opaque        q ~ hsq ~ Ct CRRulessq ~ 9psq ~ >       uq ~ A   
sq ~ Ct CRKeyq ~ Fsq ~ Ct CRValuesq ~ 9psq ~ >       uq ~ A   
sq ~ Ct Pathq ~ Fsq ~ Ct ANameq ~ Fsq ~ Ct Rulesq ~ 9psq ~ >       uq ~ A   sq ~ Cq ~ zq ~ Fsq ~ Ct Nameq ~ Fsq ~ Ct Descriptionq ~ Fsq ~ Ct AutoGenq ~ Wsq ~ Ct ReadProtq ~ Wsq ~ Ct Whileq ~ Wsq ~ Ct Nocrq ~ Wsq ~ Ct Prtyq ~ Isq ~ Ct InitUseq ~ Isq ~ Ct OnChUseq ~ Wsq ~ Ct OnChOq ~ Wpppppppppxsq ~ ?@     w      q ~ �q ~ �q ~ zq ~ ~q ~ �q ~ �q ~ �q ~ �q ~ �q ~ �q ~ �q ~ �q ~ �q ~ �q ~ �q ~ q ~ �q ~ �q ~ �q ~ �q ~ �q ~ �xq ~ z         psq ~ Ct SRefq ~ Wsq ~ Ct Aggrq ~ Wsq ~ Ct OrgAttrq ~ Fppppxsq ~ ?@     w      q ~ �q ~ �q ~ �q ~ �q ~ vq ~ uq ~ xq ~ wq ~ zq ~ yq ~ �q ~ �xt CrossReferenceRule         pppppppppxsq ~ ?@     w      q ~ qq ~ pq ~ oq ~ nxt DomainVersionCrossRefRules         psq ~ Ct OAOsq ~ 9psq ~ >       uq ~ A   
sq ~ Ct OAKq ~ Isq ~ Ct OAVsq ~ 9psq ~ >       uq ~ A   
sq ~ Ct AIDq ~ Fsq ~ Ct AIDAq ~ Fsq ~ Ct ASEq ~ Fsq ~ Ct ASEAq ~ Fppppppxsq ~ ?@     w      q ~ �q ~ �q ~ �q ~ �q ~ �q ~ �q ~ �q ~ �xt OAuthOptions         pppppppppxsq ~ ?@     w      q ~ �q ~ �q ~ �q ~ �xt DomainVersionOAuthOptions         psq ~ Ct MailInfosq ~ 9psq ~ >       uq ~ A   sq ~ Cq ~ q ~ Fsq ~ Ct INq ~ Fsq ~ Ct MHostq ~ Fsq ~ Ct MUserq ~ Fsq ~ Ct MPswdq ~ Fsq ~ Ct MProtq ~ Isq ~ Ct MPortq ~ Isq ~ Ct MCIq ~ Isq ~ Ct MSSq ~ Wsq ~ Ct SSLq ~ Wsq ~ Ct TLSq ~ Wpppppppppxsq ~ ?@     w      q ~ �q ~ �q ~ �q ~ �q ~ �q ~ �q ~ �q ~ �q ~ �q ~ �q ~ �q ~ �q ~ �q ~ �q ~ q ~ �q ~ �q ~ �q ~ �q ~ �q ~ �q ~ �xt IncomingEmailInfo         psq ~ Ct LINFsq ~ 9psq ~ >       	uq ~ A   
sq ~ Cq ~ q ~ Fsq ~ Ct LCIsq ~ 9psq ~ >       uq ~ A   
sq ~ Ct FLANq ~ Fsq ~ Ct FONq ~ Fsq ~ Ct RFANq ~ Fsq ~ Ct SUONq ~ Fppppppxsq ~ ?@     w      q ~ �q ~ �q ~ �q ~ �q ~ �q ~ �q ~ �q ~ �xt LDAPCorrespondenceInfo         psq ~ Ct AOSLq ~ Wsq ~ Ct CINFq ~ Wsq ~ Ct LATq ~ Isq ~ Ct LFORq ~ Isq ~ Ct FBsq ~ 9psq ~ >       uq ~ A   
sq ~ Ct MPsq ~ 9psq ~ >       uq ~ A   
sq ~ Ct OFq ~ Fsq ~ Ct UAq ~ Fsq ~ Ct PRq ~ Wpppppppxsq ~ ?@     w      q ~ �q ~ �q ~ �q ~ �q ~ �q ~ �xt OAuthMapping         psq ~ Ct UOq ~ Fsq ~ Ct CAq ~ Wpppppppxsq ~ ?@     w      q ~q ~q ~q ~q ~ �q ~ �xt OAuthLoginOptions         psq ~ Ct GGLq ~ �sq ~ Ct TWq ~ �pxsq ~ ?@     w      	q ~ �q ~ �q ~ �q ~ �q ~ �q ~ �q ~ �q ~ �q ~ �q ~ �q ~q ~q ~ q ~ �q ~ �q ~ �q ~
q ~	xt 	LoginInfo         psq ~ Ct DBSsq ~ 9psq ~ >       uq ~ A   
sq ~ Cq ~ q ~ Fsq ~ Ct DBq ~ Isq ~ Ct SQLsq ~ 9psq ~ >       uq ~ A   
sq ~ Ct STMTq ~ Fpppppppppxsq ~ ?@     w      q ~q ~xt DatabaseScript_Statement         ppppppppxsq ~ ?@     w      q ~q ~q ~q ~q ~ q ~xt DatabaseScript         psq ~ Cq ~ q ~ Wsq ~ Cq ~ )q ~ Wsq ~ Cq ~ 'q ~ Wsq ~ Cq ~ #q ~ Wsq ~ Cq ~ q ~ Wpppppppxsq ~ ?@     #w   /   !q ~ q ~ [q ~ 
q ~ Hq ~ q ~$q ~ �q ~ �q ~ Zq ~ Yq ~ Uq ~ Tq ~ q ~ Eq ~ q ~ aq ~q ~q ~ q ~ Oq ~ q ~ `q ~ q ~ q ~ q ~ Vq ~ q ~ Rq ~ Mq ~ Lq ~ q ~ fq ~ !q ~ \q ~ #q ~#q ~ %q ~ Kq ~ 'q ~"q ~ +q ~ Pq ~ -q ~ _q ~ )q ~!q ~ �q ~ �q ~ �q ~ �q ~ /q ~ Nq ~ 1q ~ Qq ~ 3q ~ ]q ~ 5q ~ Sq ~ jq ~ iq ~ eq ~ dq ~ 7q ~ ^q ~ cq ~ bxt DomainVersionImpl         p